MACRO DFFAR_1X ;
CLASS CORE ;
FOREIGN DFFAR_1X 0.0 0.0 ;
ORIGIN 0.0 162.0;
SIZE 648.0 BY 0.0;
SYMMETRY X Y ;
SITE UNIT ;

PIN CLK ;
DIRECTION INPUT ;
PORT
LAYER M1 ;
RECT 17.5 8.5 18.5 9.5
END
END CLK ;

PIN DATA ;
DIRECTION INPUT ;
PORT
LAYER M1 ;
RECT 125.5 8.5 126.5 9.5
END
END DATA ;

PIN NRST ;
DIRECTION INPUT ;
PORT
LAYER M1 ;
RECT 305.5 8.5 306.5 9.5
END
END NRST ;

PIN OUT ;
DIRECTION INPUT ;
PORT
LAYER M1 ;
RECT 617.5 104.5 618.5 105.5
END
END OUT ;

PIN VDD ;
USE GROUND ;
PORT
LAYER M1 ;
RECT 41.5 152.5 42.5 153.5 ;
RECT 89.5 152.5 90.5 153.5 ;
RECT 113.5 152.5 114.5 153.5 ;
RECT 257.5 152.5 258.5 153.5 ;
RECT 329.5 152.5 330.5 153.5 ;
RECT 341.5 152.5 342.5 153.5 ;
RECT 485.5 152.5 486.5 153.5 ;
RECT 473.5 152.5 474.5 153.5 ;
RECT 581.5 152.5 582.5 153.5 ;
RECT -0.5 140.5 0.5 141.5 ;
RECT 629.5 152.5 630.5 153.5 ;
END
END VDD

PIN VSS ;
USE GROUND ;
PORT
LAYER M1 ;
RECT 3.0 18.0 9.0 24.0 ;
RECT 39.0 18.0 45.0 24.0 ;
RECT 87.0 18.0 93.0 24.0 ;
RECT 111.0 18.0 117.0 24.0 ;
RECT 255.0 18.0 261.0 24.0 ;
RECT 339.0 18.0 345.0 24.0 ;
RECT 483.0 18.0 489.0 24.0 ;
RECT 471.0 18.0 477.0 24.0 ;
RECT 507.0 18.0 513.0 24.0 ;
RECT 579.0 18.0 585.0 24.0 ;
RECT 627.0 18.0 633.0 24.0 ;
RECT -3.0 18.0 3.0 24.0 ;
END
END VSS

OBS 
LAYER M1 ;
RECT 15.0 102.0 21.0 108.0
RECT 15.0 54.0 21.0 60.0
RECT 3.0 126.0 9.0 132.0
RECT 51.0 54.0 57.0 60.0
RECT 51.0 126.0 57.0 132.0
RECT 63.0 54.0 69.0 60.0
RECT 75.0 54.0 81.0 60.0
RECT 63.0 90.0 69.0 96.0
RECT 75.0 102.0 81.0 108.0
RECT 171.0 102.0 177.0 108.0
RECT 159.0 102.0 165.0 108.0
RECT 123.0 54.0 129.0 60.0
RECT 123.0 102.0 129.0 108.0
RECT 135.0 126.0 141.0 132.0
RECT 135.0 54.0 141.0 60.0
RECT 159.0 54.0 165.0 60.0
RECT 183.0 102.0 189.0 108.0
RECT 183.0 90.0 189.0 96.0
RECT 183.0 54.0 189.0 60.0
RECT 183.0 54.0 189.0 60.0
RECT 195.0 66.0 201.0 72.0
RECT 231.0 102.0 237.0 108.0
RECT 267.0 102.0 273.0 108.0
RECT 219.0 114.0 225.0 120.0
RECT 219.0 114.0 225.0 120.0
RECT 279.0 114.0 285.0 120.0
RECT 195.0 126.0 201.0 132.0
RECT 267.0 66.0 273.0 72.0
RECT 303.0 54.0 309.0 60.0
RECT 303.0 102.0 309.0 108.0
RECT 207.0 90.0 213.0 96.0
RECT 207.0 54.0 213.0 60.0
RECT 195.0 42.0 201.0 48.0
RECT 291.0 102.0 297.0 108.0
RECT 279.0 90.0 285.0 96.0
RECT 279.0 54.0 285.0 60.0
RECT 231.0 30.0 237.0 36.0
RECT 231.0 54.0 237.0 60.0
RECT 291.0 54.0 297.0 60.0
RECT 363.0 102.0 369.0 108.0
RECT 351.0 90.0 357.0 96.0
RECT 351.0 54.0 357.0 60.0
RECT 363.0 54.0 369.0 60.0
RECT 75.0 78.0 81.0 84.0
RECT 375.0 102.0 381.0 108.0
RECT 387.0 54.0 393.0 60.0
RECT 3.0 126.0 9.0 132.0
RECT 399.0 102.0 405.0 108.0
RECT 399.0 90.0 405.0 96.0
RECT 399.0 54.0 405.0 60.0
RECT 399.0 54.0 405.0 60.0
RECT 411.0 126.0 417.0 132.0
RECT 423.0 90.0 429.0 96.0
RECT 423.0 54.0 429.0 60.0
RECT 291.0 66.0 297.0 72.0
RECT 291.0 66.0 297.0 72.0
RECT 351.0 66.0 357.0 72.0
RECT 519.0 54.0 525.0 60.0
RECT 555.0 54.0 561.0 60.0
RECT 555.0 102.0 561.0 108.0
RECT 591.0 102.0 597.0 108.0
RECT 519.0 102.0 525.0 108.0
RECT 411.0 42.0 417.0 48.0
RECT 375.0 42.0 381.0 48.0
RECT 387.0 126.0 393.0 132.0
RECT 303.0 30.0 309.0 36.0
RECT 195.0 66.0 201.0 72.0
RECT 447.0 78.0 453.0 84.0
RECT 591.0 90.0 597.0 96.0
RECT 447.0 102.0 453.0 108.0
RECT 531.0 54.0 537.0 60.0
RECT 531.0 90.0 537.0 96.0
RECT 543.0 54.0 549.0 60.0
RECT 591.0 78.0 597.0 84.0
RECT 411.0 66.0 417.0 72.0
RECT 411.0 66.0 417.0 72.0
RECT 555.0 66.0 561.0 72.0
RECT 435.0 54.0 441.0 60.0
END

END  DFFAR_1X
